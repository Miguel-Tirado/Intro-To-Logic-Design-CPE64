module comparatorv2_tb();
	reg a0,a1,a2,b0,b1,b2;
	wire G,E,L;
	
	comparatorv2 uut (.a0(a0), .a1(a1), .a2(a2), .b0(b0), .b1(b1), .b2(b2), .G(G), .E(E), .L(L));
	
	initial begin 
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b0;b2 = 1'b0; b1 = 1'b0; b0 = 1'b0; //0
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b0;b2 = 1'b0; b1 = 1'b0; b0 = 1'b1; //1
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b0;b2 = 1'b0; b1 = 1'b1; b0 = 1'b0; //2
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b0;b2 = 1'b0; b1 = 1'b1; b0 = 1'b1; //3
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b0;b2 = 1'b1; b1 = 1'b0; b0 = 1'b0; //4
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b0;b2 = 1'b1; b1 = 1'b0; b0 = 1'b1; //5jj
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b0;b2 = 1'b1; b1 = 1'b1; b0 = 1'b0; //6
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b0;b2 = 1'b1; b1 = 1'b1; b0 = 1'b1; //7
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b1;b2 = 1'b0; b1 = 1'b0; b0 = 1'b0; //8
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b1;b2 = 1'b0; b1 = 1'b0; b0 = 1'b1; //9
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b1;b2 = 1'b0; b1 = 1'b1; b0 = 1'b0; //10
	#20
	a2 = 1'b0;a1 = 1'b0;a0 = 1'b1;b2 = 1'b0; b1 = 1'b1; b0 = 1'b1; //11
	#20;
	
 end 
endmodule 