module notgate(in1,out);
	input in1;
	output out;
	
	wire in1, out;
	
	not g1(out,in1);
	
endmodule 